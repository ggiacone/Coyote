
 //
	// USER LOGIC
//

ternaryGEMMOP inst_user_logic_GEMM (

        .axi_ctrl_awvalid(axi_ctrl.awvalid),
        .axi_ctrl_awready(axi_ctrl.awready),
        .axi_ctrl_awaddr(axi_ctrl.awaddr),
        .axi_ctrl_awprot(),
        .axi_ctrl_wvalid(axi_ctrl.wvalid),
        .axi_ctrl_wready(axi_ctrl.wready),
        .axi_ctrl_wdata(axi_ctrl.wdata),
        .axi_ctrl_wstrb(axi_ctrl.wstrb),
        .axi_ctrl_arvalid(axi_ctrl.arvalid),
        .axi_ctrl_arready(axi_ctrl.arready),
        .axi_ctrl_araddr(axi_ctrl.araddr),
        .axi_ctrl_arprot(),
        .axi_ctrl_rvalid(axi_ctrl.rvalid),
        .axi_ctrl_rready(axi_ctrl.ready),
        .axi_ctrl_rdata(axi_ctrl.rdata),
        .axi_ctrl_rresp(axi_ctrl.rresp),
        .axi_ctrl_bvalid(axi_ctrl.bvalid),
        .axi_ctrl_bready(axi_ctrl.bready),
        .axi_ctrl_bresp(axi_ctrl.bresp),

        .hostd_bpss_rd_req_data(sq_rd.data),
        .hostd_bpss_rd_req_valid(sq_rd.valid),
        .hostd_bpss_rd_req_ready(sq_rd.ready),
        .hostd_bpss_wr_req_data(sq_wr.data),
        .hostd_bpss_wr_req_valid(sq_wr.valid),
        .hostd_bpss_wr_req_ready(sq_wr.ready),
        .hostd_bpss_rd_done_data(cq_rd.data),
        .hostd_bpss_rd_done_valid(cq_rd.valid),
        .hostd_bpss_rd_done_ready(),
        .hostd_bpss_wr_done_data(cq_wr.data),
        .hostd_bpss_wr_done_valid(cq_wr.valid),
        .hostd_bpss_wr_done_ready(),

        .hostd_axis_host_sink_tdata(axis_host_recv[0].tdata),
        .hostd_axis_host_sink_tkeep(axis_host_recv[0].tkeep),
        .hostd_axis_host_sink_tdest(axis_host_recv[0].tid),
        .hostd_axis_host_sink_tlast(axis_host_recv[0].tlast),
        .hostd_axis_host_sink_tvalid(axis_host_recv[0].tvalid),
        .hostd_axis_host_sink_tready(axis_host_recv[0].tready),
        .hostd_axis_host_src_tdata(axis_host_send[0].tdata),
        .hostd_axis_host_src_tkeep(axis_host_send[0].tkeep),
        .hostd_axis_host_src_tdest(axis_host_send[0].tid),
        .hostd_axis_host_src_tlast(axis_host_send[0].tlast),
        .hostd_axis_host_src_tvalid(axis_host_send[0].tvalid),
        .hostd_axis_host_src_tready(axis_host_send[0].tready),
# waiting for shien
            .axi_mem_0_awvalid(axi_mem_0_awvalid),
            .axi_mem_0_awready(axi_mem_0_awready),
            .axi_mem_0_awaddr(axi_mem_0_awaddr),
            .axi_mem_0_awid(axi_mem_0_awid),
            .axi_mem_0_awlen(axi_mem_0_awlen),
            .axi_mem_0_awsize(axi_mem_0_awsize),
            .axi_mem_0_awburst(axi_mem_0_awburst),

            .axi_mem_0_wvalid(axi_mem_0_wvalid),
            .axi_mem_0_wready(axi_mem_0_wready),
            .axi_mem_0_wdata(axi_mem_0_wdata),
            .axi_mem_0_wstrb(axi_mem_0_wstrb),
            .axi_mem_0_wlast(axi_mem_0_wlast),
            .axi_mem_0_bvalid(axi_mem_0_bvalid),
            .axi_mem_0_bready(axi_mem_0_bready),
            .axi_mem_0_bid(axi_mem_0_bid),
            .axi_mem_0_bresp(axi_mem_0_bresp),

            .axi_mem_0_arvalid(axi_mem_0_arvalid),
            .axi_mem_0_arready(axi_mem_0_arready),
            .axi_mem_0_araddr(axi_mem_0_araddr),
            .axi_mem_0_arid(axi_mem_0_arid),
            .axi_mem_0_arlen(axi_mem_0_arlen),
            .axi_mem_0_arsize(axi_mem_0_arsize),
            .axi_mem_0_arburst(axi_mem_0_arburst),

            .axi_mem_0_rvalid(axi_mem_0_rvalid),
            .axi_mem_0_rready(axi_mem_0_rready),
            .axi_mem_0_rdata(axi_mem_0_rdata),
            .axi_mem_0_rid(axi_mem_0_rid),
            .axi_mem_0_rresp(axi_mem_0_rresp),
            .axi_mem_0_rlast(axi_mem_0_rlast),

            .axi_mem_1_awvalid(axi_mem_1_awvalid),
            .axi_mem_1_awready(axi_mem_1_awready),
            .axi_mem_1_awaddr(axi_mem_1_awaddr),
            .axi_mem_1_awid(axi_mem_1_awid),
            .axi_mem_1_awlen(axi_mem_1_awlen),
            .axi_mem_1_awsize(axi_mem_1_awsize),
            .axi_mem_1_awburst(axi_mem_1_awburst),

            .axi_mem_1_wvalid(axi_mem_1_wvalid),
            .axi_mem_1_wready(axi_mem_1_wready),
            .axi_mem_1_wdata(axi_mem_1_wdata),
            .axi_mem_1_wstrb(axi_mem_1_wstrb),
            .axi_mem_1_wlast(axi_mem_1_wlast),
            .axi_mem_1_bvalid(axi_mem_1_bvalid),
            .axi_mem_1_bready(axi_mem_1_bready),
            .axi_mem_1_bid(axi_mem_1_bid),
            .axi_mem_1_bresp(axi_mem_1_bresp),

            .axi_mem_1_arvalid(axi_mem_1_arvalid),
            .axi_mem_1_arready(axi_mem_1_arready),
            .axi_mem_1_araddr(axi_mem_1_araddr),
            .axi_mem_1_arid(axi_mem_1_arid),
            .axi_mem_1_arlen(axi_mem_1_arlen),
            .axi_mem_1_arsize(axi_mem_1_arsize),
            .axi_mem_1_arburst(axi_mem_1_arburst),

            .axi_mem_1_rvalid(exiaxi_mem_1_rvalid),
            .axi_mem_1_rready(axi_mem_1_rready),
            .axi_mem_1_rdata(axi_mem_1_rdata),
            .axi_mem_1_rid(axi_mem_1_rid),
            .axi_mem_1_rresp(axi_mem_1_rresp),
            .axi_mem_1_rlast(axi_mem_1_rlast),

        .resetn(aresetn),
        .clk(aclk)
	);
